module tb_top_MBE();
	parameter int unsigned NBIT = 23;
	parameter int unsigned NBLOCK = 9;

	logic [NBIT:0] i_X, i_Y;
	logic [47:0] o_P;

	top_MBE_R8 #(
		.NBIT_MANTISSA(NBIT),
		.NBLOCK(NBLOCK)
	)  C_MBE (
		.X(i_X),
		.Y(i_Y),
		.P(o_P)
	);

	initial
	begin
		#10
		i_X = 24'b111100000000000000001110;		//      full-->111100000000000000001110=15728654
		i_Y = 24'b100000001010110000010100;		//      full-->100000001010110000010100=8432660
												// 132,634,391,439,640
		#10
		i_X = 24'b111100000000000000001110;		//       full-->111100000000000000001110=15728654
		i_Y = 24'b100000000000000110010100;		//       full-->100000000000000110010100=8389012
												//   131,947,867,149,848

		#10
		i_X = 24'b111111111111111111111111;		//       full-->111111111111111111111111=16777215
        i_Y = 24'b111111111111111111111111;		//       full-->111111111111111111111111=16777215  
												// 281,474,943,156,225
		#10
		i_X = 24'b111110010111111001010100;      //      full-->111110010111111001010100=16350804
	    i_Y = 24'd0;                            //       full-->100000000000000000000000=8388608
                                                //  137,160,485,240,832     
	    #10
	    i_X = $random;                       //verify in report
	    i_Y = $random;
	    #10
	    i_X = $random;
	    i_Y = $random;

	     #10
	    i_X = $random;
	    i_Y = $random;

	     #10
	    i_X = $random;
	    i_Y = $random;

	     #10
	    i_X = $random;
	    i_Y = $random;

	    
       

	end
endmodule